module toInst
(
  parameter width_sdajdads = 25,
  parameter width2_asdf = 30
)
(
  input [2-1:0] aasdasd,
  input [2-1:0] bdasdasf,
  output reg [width2_asdf-1:0] cfafafafasf
);
endmodule;
