always_ff @( clock ) begin : blockName
    case
        
    endcase
end
