always_ff @( clock ) begin : blockName
    case
        
    endcase
end
always_comb begin : tea
    a = 
end
// a is a variable
reg k; // after comment

always_comb begin
    k = 33;
end

toInst u_toInst(
	.a(a),
    .b(b),
    .c(c)
);

toInst 
#(
    .width(width),
    .width2(width2)
)
u_toInst(
	.a(a),
    .b(b),
    .c(c)
);

mod_name instance_name (.*);
toInst 
#(
    .width_sdajdads (width_sdajdads ),
    .width2_asdf    (width2_asdf    )
)
u_toInst(
	.aasdasd     (aasdasd     ),
    .bdasdasf    (bdasdasf    ),
    .cfafafafasf (cfafafafasf )
);

/*
dasdas
dasda
*/
// sdas
  reg aa=15; 
  reg aaa= 33; 

  wire [13:fd0] aa; 
  wire [hkjghj-45:  0] bb; 
  wire [fsdfsfs-255:  0] vv; //sdfsfs
  reg  [12:ghjds+1] dd [35:15];//wire reg a = fdfds; 

  assign a={dd[15][24:0],dd[14][64:9]} ; 
  assign b=35848+fsfsf; 


always_comb begin
  a= 15; 
  addfdf = 33 ; 
      fff= 15 + gfdg; 
  dsfs[7487:46]=fsdfs[fsdf]+fsdfs+fsfsd;
end

always_ff(@posedge clk)begin
  {a[65:314],b[fdsf:577]}<= 57; 
  c[15:0]    <= df; 
  fsdf <= df+fsdfs; 
  if(fsdfsd)begin
    dfdsf<= {df+fsdfsd, sfds[das:dasdas}; 
  end
  else begin
    dfsdf <=fdfdsfsfs; 
    fdsfds<=dsfsdfs  ; 
  end
end

aa
toInst 
#(
    .width_sdajdads (width_sdajdads ),
    .width2_asdf    (width2_asdf    )
)
u_toInst(
	.aasdasd     (aasdasd     ),
    .bdasdasf    (bdasdasf    ),
    .cfafafafasf (cfafafafasf )
);

